
module CELL_BLOCK #(parameter DATA_WIDTH = 14, OUTPUT_WIDTH = 14) (
    input wire clk, rst,
    input wire store_enable,
    input wire [DATA_WIDTH-1:0] i,
    input wire [DATA_WIDTH-1:0] f,
    input wire [DATA_WIDTH-1:0] c,
    
    output reg [DATA_WIDTH-1:0] cell_state
);

reg [DATA_WIDTH-1:0] cell_state_old;

wire [2*DATA_WIDTH-1:0] mult1;
wire [2*DATA_WIDTH-1:0] mult2;
wire [2*DATA_WIDTH-1:0] cell_state_large;
wire [1*DATA_WIDTH-1:0] cell_state_small;

WallaceTreeMul MULT1(f, cell_state_old, mult1);
WallaceTreeMul MULT2(i, c,              mult2);

Kogge_Stone_ADDER_28 ADD1(mult1, mult2, 1'b0, cell_state_large);
Kogge_Stone_ADDER_14 ADD1_R(cell_state_large[23:10], 14'b0_000_0000000000, cell_state_large[9], cell_state_small);

always @(*) begin
    cell_state = cell_state_small;
end

always @(posedge clk or negedge rst) begin
    if(!rst) begin
        cell_state_old <= 14'b0_000_0000000000;
    end
    else begin
        if(store_enable) begin
            cell_state_old <= cell_state_small;
        end
    end
end

endmodule


/////////////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////


module HIDDEN_BLOCK #(parameter DATA_WIDTH = 14, OUTPUT_WIDTH = 14) (
    input wire clk, rst,
    input wire store_hidden_enable,
    input wire [DATA_WIDTH-1:0] cell_state,
    input wire [DATA_WIDTH-1:0] o,

    output reg [DATA_WIDTH-1:0] hidden_state
);

wire [DATA_WIDTH-1:0] tanh_out;
wire [2*DATA_WIDTH-1:0] mult1;
wire [DATA_WIDTH-1:0] hidden_state_reg;
reg [DATA_WIDTH-1:0] o_reg;

always @(posedge clk or negedge rst) begin
    if(!rst) begin
        o_reg <= 14'b0_000_0000000000;
    end
    else begin
        o_reg <= o;
    end
end

Tanh_TOP_H TANH(clk, rst, cell_state, tanh_out);
WallaceTreeMul MULT1(tanh_out, o_reg, mult1);

Kogge_Stone_ADDER_14 ADD1_R(mult1[23:10], 14'b0_000_0000000000, mult1[9], hidden_state_reg);

always @(posedge clk or negedge rst) begin
    if(!rst) begin
        hidden_state <= 14'b0_000_0000000000;
    end
    else begin
        if(store_hidden_enable == 1'b1) begin
            hidden_state <= hidden_state_reg;
        end
    end
end
    
endmodule


//////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////////////




module CELL_HIDDEN_BLOCK #(parameter DATA_WIDTH = 14, OUTPUT_WIDTH = 14) (
    input wire clk, rst,
    input wire store_enable,
    input wire store_hidden_enable,
    input wire [DATA_WIDTH-1:0] i,
    input wire [DATA_WIDTH-1:0] f,
    input wire [DATA_WIDTH-1:0] c,
    input wire [DATA_WIDTH-1:0] o,

    output wire [DATA_WIDTH-1:0] hidden_state
);

wire [DATA_WIDTH-1:0] cell_state;
CELL_BLOCK CSB (clk, rst, store_enable, i, f, c, cell_state);
HIDDEN_BLOCK HSB (clk, rst, store_hidden_enable, cell_state, o, hidden_state);

endmodule